library verilog;
use verilog.vl_types.all;
entity test_cla4bit is
end test_cla4bit;
